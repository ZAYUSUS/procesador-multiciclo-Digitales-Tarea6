module MemDataReg (
    input [31:0] inst,
    output  [63:0] Mem_data_reg
);
    assign Mem_data_reg=0;
endmodule